----------------------------------------------------------------------------------
-- This file has been mechanically generated
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OffsetTable is
	port(
		addr_i	: in std_logic_vector(9 downto 0);
		data_o	: out std_logic_vector(19 downto 0)
	);
end entity;

architecture procedural of OffsetTable is
begin
	P_look_up : process(addr_i)
	begin
		case addr_i is
			when "1000000000" => data_o <= "11111111000000000000";
			when "1000000001" => data_o <= "11111111000000000000";
			when "1000000010" => data_o <= "11111111000000000000";
			when "1000000011" => data_o <= "11111111000000000000";
			when "1000000100" => data_o <= "11111111000000000000";
			when "1000000101" => data_o <= "11111111000000000000";
			when "1000000110" => data_o <= "11111111000000000000";
			when "1000000111" => data_o <= "11111111000000000000";
			when "1000001000" => data_o <= "11111111000000000000";
			when "1000001001" => data_o <= "11111111000000000000";
			when "1000001010" => data_o <= "11111111000000000000";
			when "1000001011" => data_o <= "11111111000000000000";
			when "1000001100" => data_o <= "11111111000000000000";
			when "1000001101" => data_o <= "11111111000000000000";
			when "1000001110" => data_o <= "11111111000000000000";
			when "1000001111" => data_o <= "11111111000000000000";
			when "1000010000" => data_o <= "11111111000000000000";
			when "1000010001" => data_o <= "11111111000000000000";
			when "1000010010" => data_o <= "11111111000000000000";
			when "1000010011" => data_o <= "11111111000000000000";
			when "1000010100" => data_o <= "11111111000000000000";
			when "1000010101" => data_o <= "11111111000000000000";
			when "1000010110" => data_o <= "11111111000000000000";
			when "1000010111" => data_o <= "11111111000000000000";
			when "1000011000" => data_o <= "11111111000000000000";
			when "1000011001" => data_o <= "11111111000000000000";
			when "1000011010" => data_o <= "11111111000000000000";
			when "1000011011" => data_o <= "11111111000000000000";
			when "1000011100" => data_o <= "11111111000000000000";
			when "1000011101" => data_o <= "11111111000000000000";
			when "1000011110" => data_o <= "11111111000000000000";
			when "1000011111" => data_o <= "11111111000000000000";
			when "1000100000" => data_o <= "11111111000000000000";
			when "1000100001" => data_o <= "11111111000000000000";
			when "1000100010" => data_o <= "11111111000000000000";
			when "1000100011" => data_o <= "11111111000000000000";
			when "1000100100" => data_o <= "11111111000000000000";
			when "1000100101" => data_o <= "11111111000000000000";
			when "1000100110" => data_o <= "11111111000000000000";
			when "1000100111" => data_o <= "11111111000000000000";
			when "1000101000" => data_o <= "11111111000000000000";
			when "1000101001" => data_o <= "11111111000000000000";
			when "1000101010" => data_o <= "11111111000000000000";
			when "1000101011" => data_o <= "11111111000000000000";
			when "1000101100" => data_o <= "11111111000000000000";
			when "1000101101" => data_o <= "11111111000000000000";
			when "1000101110" => data_o <= "11111111000000000000";
			when "1000101111" => data_o <= "11111111000000000000";
			when "1000110000" => data_o <= "11111111000000000000";
			when "1000110001" => data_o <= "11111111000000000000";
			when "1000110010" => data_o <= "11111111000000000000";
			when "1000110011" => data_o <= "11111111000000000000";
			when "1000110100" => data_o <= "11111111000000000000";
			when "1000110101" => data_o <= "11111111000000000000";
			when "1000110110" => data_o <= "11111111000000000000";
			when "1000110111" => data_o <= "11111111000000000000";
			when "1000111000" => data_o <= "11111111000000000000";
			when "1000111001" => data_o <= "11111111000000000000";
			when "1000111010" => data_o <= "11111111000000000000";
			when "1000111011" => data_o <= "11111111000000000000";
			when "1000111100" => data_o <= "11111111000000000000";
			when "1000111101" => data_o <= "11111111000000000000";
			when "1000111110" => data_o <= "11111111000000000000";
			when "1000111111" => data_o <= "11111111000000000000";
			when "1001000000" => data_o <= "11111111000000000000";
			when "1001000001" => data_o <= "11111111000000000000";
			when "1001000010" => data_o <= "11111111000000000000";
			when "1001000011" => data_o <= "11111111000000000000";
			when "1001000100" => data_o <= "11111111000000000000";
			when "1001000101" => data_o <= "11111111000000000000";
			when "1001000110" => data_o <= "11111111000000000000";
			when "1001000111" => data_o <= "11111111000000000000";
			when "1001001000" => data_o <= "11111111000000000000";
			when "1001001001" => data_o <= "11111111000000000000";
			when "1001001010" => data_o <= "11111111000000000000";
			when "1001001011" => data_o <= "11111111000000000000";
			when "1001001100" => data_o <= "11111111000000000000";
			when "1001001101" => data_o <= "11111111000000000000";
			when "1001001110" => data_o <= "11111111000000000000";
			when "1001001111" => data_o <= "11111111000000000000";
			when "1001010000" => data_o <= "11111111000000000000";
			when "1001010001" => data_o <= "11111111000000000000";
			when "1001010010" => data_o <= "11111111000000000000";
			when "1001010011" => data_o <= "11111111000000000000";
			when "1001010100" => data_o <= "11111111000000000000";
			when "1001010101" => data_o <= "11111111000000000000";
			when "1001010110" => data_o <= "11111111000000000000";
			when "1001010111" => data_o <= "11111111000000000000";
			when "1001011000" => data_o <= "11111111000000000000";
			when "1001011001" => data_o <= "11111111000000000000";
			when "1001011010" => data_o <= "11111111000000000000";
			when "1001011011" => data_o <= "11111111000000000000";
			when "1001011100" => data_o <= "11111111000000000000";
			when "1001011101" => data_o <= "11111111000000000000";
			when "1001011110" => data_o <= "11111111000000000000";
			when "1001011111" => data_o <= "11111111000000000000";
			when "1001100000" => data_o <= "11111111000000000000";
			when "1001100001" => data_o <= "11111111000000000000";
			when "1001100010" => data_o <= "11111111000000000000";
			when "1001100011" => data_o <= "11111111000000000000";
			when "1001100100" => data_o <= "11111111000000000000";
			when "1001100101" => data_o <= "11111111000000000000";
			when "1001100110" => data_o <= "11111111000000000000";
			when "1001100111" => data_o <= "11111111000000000000";
			when "1001101000" => data_o <= "11111111000000000000";
			when "1001101001" => data_o <= "11111111000000000000";
			when "1001101010" => data_o <= "11111111000000000000";
			when "1001101011" => data_o <= "11111111000000000000";
			when "1001101100" => data_o <= "11111111000000000000";
			when "1001101101" => data_o <= "11111111000000000000";
			when "1001101110" => data_o <= "11111111000000000000";
			when "1001101111" => data_o <= "11111111000000000000";
			when "1001110000" => data_o <= "11111111000000000000";
			when "1001110001" => data_o <= "11111111000000000000";
			when "1001110010" => data_o <= "11111111000000000000";
			when "1001110011" => data_o <= "11111111000000000000";
			when "1001110100" => data_o <= "11111111000000000000";
			when "1001110101" => data_o <= "11111111000000000000";
			when "1001110110" => data_o <= "11111111000000000000";
			when "1001110111" => data_o <= "11111111000000000000";
			when "1001111000" => data_o <= "11111111000000000000";
			when "1001111001" => data_o <= "11111111000000000000";
			when "1001111010" => data_o <= "11111111000000000000";
			when "1001111011" => data_o <= "11111111000000000000";
			when "1001111100" => data_o <= "11111111000000000000";
			when "1001111101" => data_o <= "11111111000000000000";
			when "1001111110" => data_o <= "11111111000000000000";
			when "1001111111" => data_o <= "11111111000000000000";
			when "1010000000" => data_o <= "11111111000000000000";
			when "1010000001" => data_o <= "11111111000000000000";
			when "1010000010" => data_o <= "11111111000000000000";
			when "1010000011" => data_o <= "11111111000000000000";
			when "1010000100" => data_o <= "11111111000000000000";
			when "1010000101" => data_o <= "11111111000000000000";
			when "1010000110" => data_o <= "11111111000000000000";
			when "1010000111" => data_o <= "11111111000000000000";
			when "1010001000" => data_o <= "11111111000000000000";
			when "1010001001" => data_o <= "11111111000000000000";
			when "1010001010" => data_o <= "11111111000000000000";
			when "1010001011" => data_o <= "11111111000000000000";
			when "1010001100" => data_o <= "11111111000000000000";
			when "1010001101" => data_o <= "11111111000000000000";
			when "1010001110" => data_o <= "11111111000000000000";
			when "1010001111" => data_o <= "11111111000000000000";
			when "1010010000" => data_o <= "11111111000000000000";
			when "1010010001" => data_o <= "11111111000000000000";
			when "1010010010" => data_o <= "11111111000000000000";
			when "1010010011" => data_o <= "11111111000000000000";
			when "1010010100" => data_o <= "11111111000000000000";
			when "1010010101" => data_o <= "11111111000000000000";
			when "1010010110" => data_o <= "11111111000000000000";
			when "1010010111" => data_o <= "11111111000000000000";
			when "1010011000" => data_o <= "11111111000000000000";
			when "1010011001" => data_o <= "11111111000000000000";
			when "1010011010" => data_o <= "11111111000000000000";
			when "1010011011" => data_o <= "11111111000000000000";
			when "1010011100" => data_o <= "11111111000000000000";
			when "1010011101" => data_o <= "11111111000000000000";
			when "1010011110" => data_o <= "11111111000000000000";
			when "1010011111" => data_o <= "11111111000000000000";
			when "1010100000" => data_o <= "11111111000000000000";
			when "1010100001" => data_o <= "11111111000000000000";
			when "1010100010" => data_o <= "11111111000000000000";
			when "1010100011" => data_o <= "11111111000000000000";
			when "1010100100" => data_o <= "11111111000000000000";
			when "1010100101" => data_o <= "11111111000000000000";
			when "1010100110" => data_o <= "11111111000000000000";
			when "1010100111" => data_o <= "11111111000000000000";
			when "1010101000" => data_o <= "11111111000000000000";
			when "1010101001" => data_o <= "11111111000000000000";
			when "1010101010" => data_o <= "11111111000000000000";
			when "1010101011" => data_o <= "11111111000000000000";
			when "1010101100" => data_o <= "11111111000000000000";
			when "1010101101" => data_o <= "11111111000000000000";
			when "1010101110" => data_o <= "11111111000000000000";
			when "1010101111" => data_o <= "11111111000000000000";
			when "1010110000" => data_o <= "11111111000000000000";
			when "1010110001" => data_o <= "11111111000000000000";
			when "1010110010" => data_o <= "11111111000000000000";
			when "1010110011" => data_o <= "11111111000000000000";
			when "1010110100" => data_o <= "11111111000000000000";
			when "1010110101" => data_o <= "11111111000000000000";
			when "1010110110" => data_o <= "11111111000000000000";
			when "1010110111" => data_o <= "11111111000000000000";
			when "1010111000" => data_o <= "11111111000000000000";
			when "1010111001" => data_o <= "11111111000000000000";
			when "1010111010" => data_o <= "11111111000000000000";
			when "1010111011" => data_o <= "11111111000000000000";
			when "1010111100" => data_o <= "11111111000000000000";
			when "1010111101" => data_o <= "11111111000000000000";
			when "1010111110" => data_o <= "11111111000000000000";
			when "1010111111" => data_o <= "11111111000000000000";
			when "1011000000" => data_o <= "11111111000000000000";
			when "1011000001" => data_o <= "11111111000000000000";
			when "1011000010" => data_o <= "11111111000000000000";
			when "1011000011" => data_o <= "11111111000000000000";
			when "1011000100" => data_o <= "11111111000000000000";
			when "1011000101" => data_o <= "11111111000000000000";
			when "1011000110" => data_o <= "11111111000000000000";
			when "1011000111" => data_o <= "11111111000000000000";
			when "1011001000" => data_o <= "11111111000000000000";
			when "1011001001" => data_o <= "11111111000000000000";
			when "1011001010" => data_o <= "11111111000000000000";
			when "1011001011" => data_o <= "11111111000000000000";
			when "1011001100" => data_o <= "11111111000000000000";
			when "1011001101" => data_o <= "11111111000000000000";
			when "1011001110" => data_o <= "11111111000000000000";
			when "1011001111" => data_o <= "11111111000000000000";
			when "1011010000" => data_o <= "11111111000000000000";
			when "1011010001" => data_o <= "11111111000000000000";
			when "1011010010" => data_o <= "11111111000000000000";
			when "1011010011" => data_o <= "11111111000000000000";
			when "1011010100" => data_o <= "11111111000000000000";
			when "1011010101" => data_o <= "11111111000000000000";
			when "1011010110" => data_o <= "11111111000000000000";
			when "1011010111" => data_o <= "11111111000000000000";
			when "1011011000" => data_o <= "11111111000000000000";
			when "1011011001" => data_o <= "11111111000000000000";
			when "1011011010" => data_o <= "11111111000000000000";
			when "1011011011" => data_o <= "11111111000000000000";
			when "1011011100" => data_o <= "11111111000000000000";
			when "1011011101" => data_o <= "11111111000000000000";
			when "1011011110" => data_o <= "11111111000000000000";
			when "1011011111" => data_o <= "11111111000000000000";
			when "1011100000" => data_o <= "11111111000000000000";
			when "1011100001" => data_o <= "11111111000000000000";
			when "1011100010" => data_o <= "11111111000000000000";
			when "1011100011" => data_o <= "11111111000000000000";
			when "1011100100" => data_o <= "11111111000000000000";
			when "1011100101" => data_o <= "11111111000000000000";
			when "1011100110" => data_o <= "11111111000000000000";
			when "1011100111" => data_o <= "11111111000000000000";
			when "1011101000" => data_o <= "11111111000000000000";
			when "1011101001" => data_o <= "11111111000000000000";
			when "1011101010" => data_o <= "11111111000000000000";
			when "1011101011" => data_o <= "11111111000000000000";
			when "1011101100" => data_o <= "11111111000000000000";
			when "1011101101" => data_o <= "11111111000000000000";
			when "1011101110" => data_o <= "11111111000000000000";
			when "1011101111" => data_o <= "11111111000000000000";
			when "1011110000" => data_o <= "11111111000000000000";
			when "1011110001" => data_o <= "11111111000000000000";
			when "1011110010" => data_o <= "11111111000000000000";
			when "1011110011" => data_o <= "11111111000000000000";
			when "1011110100" => data_o <= "11111111000000000000";
			when "1011110101" => data_o <= "11111111000000000000";
			when "1011110110" => data_o <= "11111111000000000000";
			when "1011110111" => data_o <= "11111111000000000000";
			when "1011111000" => data_o <= "11111111000000000000";
			when "1011111001" => data_o <= "11111111000000000000";
			when "1011111010" => data_o <= "11111111000000000000";
			when "1011111011" => data_o <= "11111111000000000000";
			when "1011111100" => data_o <= "11111111000000000000";
			when "1011111101" => data_o <= "11111111000000000000";
			when "1011111110" => data_o <= "11111111000000000000";
			when "1011111111" => data_o <= "11111111000000000000";
			when "1100000000" => data_o <= "11111111000000000000";
			when "1100000001" => data_o <= "11111111000000000000";
			when "1100000010" => data_o <= "11111111000000000000";
			when "1100000011" => data_o <= "11111111000000000000";
			when "1100000100" => data_o <= "11111111000000000000";
			when "1100000101" => data_o <= "11111111000000000000";
			when "1100000110" => data_o <= "11111111000000000000";
			when "1100000111" => data_o <= "11111111000000000000";
			when "1100001000" => data_o <= "11111111000000000000";
			when "1100001001" => data_o <= "11111111000000000000";
			when "1100001010" => data_o <= "11111111000000000000";
			when "1100001011" => data_o <= "11111111000000000000";
			when "1100001100" => data_o <= "11111111000000000000";
			when "1100001101" => data_o <= "11111111000000000000";
			when "1100001110" => data_o <= "11111111000000000000";
			when "1100001111" => data_o <= "11111111000000000000";
			when "1100010000" => data_o <= "11111111000000000000";
			when "1100010001" => data_o <= "11111111000000000000";
			when "1100010010" => data_o <= "11111111000000000000";
			when "1100010011" => data_o <= "11111111000000000000";
			when "1100010100" => data_o <= "11111111000000000000";
			when "1100010101" => data_o <= "11111111000000000000";
			when "1100010110" => data_o <= "11111111000000000000";
			when "1100010111" => data_o <= "11111111000000000000";
			when "1100011000" => data_o <= "11111111000000000000";
			when "1100011001" => data_o <= "11111111000000000000";
			when "1100011010" => data_o <= "11111111000000000000";
			when "1100011011" => data_o <= "11111111000000000000";
			when "1100011100" => data_o <= "11111111000000000000";
			when "1100011101" => data_o <= "11111111000000000000";
			when "1100011110" => data_o <= "11111111000000000000";
			when "1100011111" => data_o <= "11111111000000000000";
			when "1100100000" => data_o <= "11111111000000000000";
			when "1100100001" => data_o <= "11111111000000000000";
			when "1100100010" => data_o <= "11111111000000000000";
			when "1100100011" => data_o <= "11111111000000000000";
			when "1100100100" => data_o <= "11111111000000000000";
			when "1100100101" => data_o <= "11111111000000000000";
			when "1100100110" => data_o <= "11111111000000000000";
			when "1100100111" => data_o <= "11111111000000000000";
			when "1100101000" => data_o <= "11111111000000000000";
			when "1100101001" => data_o <= "11111111000000000000";
			when "1100101010" => data_o <= "11111111000000000000";
			when "1100101011" => data_o <= "11111111000000000000";
			when "1100101100" => data_o <= "11111111000000000000";
			when "1100101101" => data_o <= "11111111000000000000";
			when "1100101110" => data_o <= "11111111000000000000";
			when "1100101111" => data_o <= "11111111000000000000";
			when "1100110000" => data_o <= "11111111000000000000";
			when "1100110001" => data_o <= "11111111000000000000";
			when "1100110010" => data_o <= "11111111000000000000";
			when "1100110011" => data_o <= "11111111000000000000";
			when "1100110100" => data_o <= "11111111000000000000";
			when "1100110101" => data_o <= "11111111000000000000";
			when "1100110110" => data_o <= "11111111000000000000";
			when "1100110111" => data_o <= "11111111000000000000";
			when "1100111000" => data_o <= "11111111000000000000";
			when "1100111001" => data_o <= "11111111000000000000";
			when "1100111010" => data_o <= "11111111000000000000";
			when "1100111011" => data_o <= "11111111000000000000";
			when "1100111100" => data_o <= "11111111000000000000";
			when "1100111101" => data_o <= "11111111000000000000";
			when "1100111110" => data_o <= "11111111000000000000";
			when "1100111111" => data_o <= "11111111000000000000";
			when "1101000000" => data_o <= "11111111000000000000";
			when "1101000001" => data_o <= "11111111000000000000";
			when "1101000010" => data_o <= "11111111000000000000";
			when "1101000011" => data_o <= "11111111000000000000";
			when "1101000100" => data_o <= "11111111000000000000";
			when "1101000101" => data_o <= "11111111000000000000";
			when "1101000110" => data_o <= "11111111000000000000";
			when "1101000111" => data_o <= "11111111000000000000";
			when "1101001000" => data_o <= "11111111000000000000";
			when "1101001001" => data_o <= "11111111000000000000";
			when "1101001010" => data_o <= "11111111000000000000";
			when "1101001011" => data_o <= "11111111000000000000";
			when "1101001100" => data_o <= "11111111000000000000";
			when "1101001101" => data_o <= "11111111000000000000";
			when "1101001110" => data_o <= "11111111000000000000";
			when "1101001111" => data_o <= "11111111000000000000";
			when "1101010000" => data_o <= "11111111000000000000";
			when "1101010001" => data_o <= "11111111000000000000";
			when "1101010010" => data_o <= "11111111000000000000";
			when "1101010011" => data_o <= "11111111000000000000";
			when "1101010100" => data_o <= "11111111000000000000";
			when "1101010101" => data_o <= "11111111000000000000";
			when "1101010110" => data_o <= "11111111000000000000";
			when "1101010111" => data_o <= "11111111000000000000";
			when "1101011000" => data_o <= "11111111000000000000";
			when "1101011001" => data_o <= "11111111000000000000";
			when "1101011010" => data_o <= "11111111000000000000";
			when "1101011011" => data_o <= "11111111000000000000";
			when "1101011100" => data_o <= "11111111000000000000";
			when "1101011101" => data_o <= "11111111000000000000";
			when "1101011110" => data_o <= "11111111000000000000";
			when "1101011111" => data_o <= "11111111000000000000";
			when "1101100000" => data_o <= "11111111000000000000";
			when "1101100001" => data_o <= "11111111000000000000";
			when "1101100010" => data_o <= "11111111000000000000";
			when "1101100011" => data_o <= "11111111000000000000";
			when "1101100100" => data_o <= "11111111000000000000";
			when "1101100101" => data_o <= "11111111000000000000";
			when "1101100110" => data_o <= "11111111000000000000";
			when "1101100111" => data_o <= "11111111000000000000";
			when "1101101000" => data_o <= "11111111000000000000";
			when "1101101001" => data_o <= "11111111000000000000";
			when "1101101010" => data_o <= "11111111000000000000";
			when "1101101011" => data_o <= "11111111000000000000";
			when "1101101100" => data_o <= "11111111000000000000";
			when "1101101101" => data_o <= "11111111000000000000";
			when "1101101110" => data_o <= "11111111000000000000";
			when "1101101111" => data_o <= "11111111000000000000";
			when "1101110000" => data_o <= "11111111000000000000";
			when "1101110001" => data_o <= "11111111000000000000";
			when "1101110010" => data_o <= "11111111000000000000";
			when "1101110011" => data_o <= "11111111000000000000";
			when "1101110100" => data_o <= "11111111000000000000";
			when "1101110101" => data_o <= "11111111000000000000";
			when "1101110110" => data_o <= "11111111000000000000";
			when "1101110111" => data_o <= "11111111000000000000";
			when "1101111000" => data_o <= "11111111000000000000";
			when "1101111001" => data_o <= "11111111000000000000";
			when "1101111010" => data_o <= "11111111000000000000";
			when "1101111011" => data_o <= "11111111000000000000";
			when "1101111100" => data_o <= "11111111000000000000";
			when "1101111101" => data_o <= "11111111000000000000";
			when "1101111110" => data_o <= "11111111000000000000";
			when "1101111111" => data_o <= "11111111000000000000";
			when "1110000000" => data_o <= "11111111000000000000";
			when "1110000001" => data_o <= "11111111000000000000";
			when "1110000010" => data_o <= "11111111000000000000";
			when "1110000011" => data_o <= "11111111000000000000";
			when "1110000100" => data_o <= "11111111000000000000";
			when "1110000101" => data_o <= "11111111000000000000";
			when "1110000110" => data_o <= "11111111000000000000";
			when "1110000111" => data_o <= "11111111000000000000";
			when "1110001000" => data_o <= "11111111000000000000";
			when "1110001001" => data_o <= "11111111000000000000";
			when "1110001010" => data_o <= "11111111000000000000";
			when "1110001011" => data_o <= "11111111000000000000";
			when "1110001100" => data_o <= "11111111000000000000";
			when "1110001101" => data_o <= "11111111000000000000";
			when "1110001110" => data_o <= "11111111000000000000";
			when "1110001111" => data_o <= "11111111000000000000";
			when "1110010000" => data_o <= "11111111000000000000";
			when "1110010001" => data_o <= "11111111000000000000";
			when "1110010010" => data_o <= "11111111000000000000";
			when "1110010011" => data_o <= "11111111000000000000";
			when "1110010100" => data_o <= "11111111000000000000";
			when "1110010101" => data_o <= "11111111000000000000";
			when "1110010110" => data_o <= "11111111000000000000";
			when "1110010111" => data_o <= "11111111000000000000";
			when "1110011000" => data_o <= "11111111000000000000";
			when "1110011001" => data_o <= "11111111000000000000";
			when "1110011010" => data_o <= "11111111000000000000";
			when "1110011011" => data_o <= "11111111000000000000";
			when "1110011100" => data_o <= "11111111000000000000";
			when "1110011101" => data_o <= "11111111000000000000";
			when "1110011110" => data_o <= "11111111000000000000";
			when "1110011111" => data_o <= "11111111000000000000";
			when "1110100000" => data_o <= "11111111000000000000";
			when "1110100001" => data_o <= "11111111000000000000";
			when "1110100010" => data_o <= "11111111000000000000";
			when "1110100011" => data_o <= "11111111000000000000";
			when "1110100100" => data_o <= "11111111000000000000";
			when "1110100101" => data_o <= "11111111000000000000";
			when "1110100110" => data_o <= "11111111000000000000";
			when "1110100111" => data_o <= "11111111000000000000";
			when "1110101000" => data_o <= "11111111000000000000";
			when "1110101001" => data_o <= "11111111000000000000";
			when "1110101010" => data_o <= "11111111000000000000";
			when "1110101011" => data_o <= "11111111000000000000";
			when "1110101100" => data_o <= "11111111000000000000";
			when "1110101101" => data_o <= "11111111000000000000";
			when "1110101110" => data_o <= "11111111000000000000";
			when "1110101111" => data_o <= "11111111000000000000";
			when "1110110000" => data_o <= "11111111000000000000";
			when "1110110001" => data_o <= "11111111000000000000";
			when "1110110010" => data_o <= "11111111000000000000";
			when "1110110011" => data_o <= "11111111000000000000";
			when "1110110100" => data_o <= "11111111000000000000";
			when "1110110101" => data_o <= "11111111000000000000";
			when "1110110110" => data_o <= "11111111000000000001";
			when "1110110111" => data_o <= "11111111000000000001";
			when "1110111000" => data_o <= "11111111000000000001";
			when "1110111001" => data_o <= "11111111000000000001";
			when "1110111010" => data_o <= "11111111000000000001";
			when "1110111011" => data_o <= "11111111000000000001";
			when "1110111100" => data_o <= "11111111000000000001";
			when "1110111101" => data_o <= "11111111000000000001";
			when "1110111110" => data_o <= "11111111000000000001";
			when "1110111111" => data_o <= "11111111000000000001";
			when "1111000000" => data_o <= "11111111000000000001";
			when "1111000001" => data_o <= "11111111000000000001";
			when "1111000010" => data_o <= "11111111000000000001";
			when "1111000011" => data_o <= "11111111000000000001";
			when "1111000100" => data_o <= "11111111000000000001";
			when "1111000101" => data_o <= "11111111000000000001";
			when "1111000110" => data_o <= "11111111000000000001";
			when "1111000111" => data_o <= "11111111000000000001";
			when "1111001000" => data_o <= "11111111000000000001";
			when "1111001001" => data_o <= "11111111000000000001";
			when "1111001010" => data_o <= "11111111000000000001";
			when "1111001011" => data_o <= "11111111000000000001";
			when "1111001100" => data_o <= "11111111000000000001";
			when "1111001101" => data_o <= "11111111000000000001";
			when "1111001110" => data_o <= "11111111000000000001";
			when "1111001111" => data_o <= "11111111000000000001";
			when "1111010000" => data_o <= "11111111000000000001";
			when "1111010001" => data_o <= "11111111000000000001";
			when "1111010010" => data_o <= "11111111000000000001";
			when "1111010011" => data_o <= "11111111000000000001";
			when "1111010100" => data_o <= "11111111000000000001";
			when "1111010101" => data_o <= "11111111000000000001";
			when "1111010110" => data_o <= "11111111000000000001";
			when "1111010111" => data_o <= "11111111000000000001";
			when "1111011000" => data_o <= "11111111000000000001";
			when "1111011001" => data_o <= "11111111000000000001";
			when "1111011010" => data_o <= "11111111000000000001";
			when "1111011011" => data_o <= "11111111000000000001";
			when "1111011100" => data_o <= "11111111000000000001";
			when "1111011101" => data_o <= "11111111000000000001";
			when "1111011110" => data_o <= "11111111000000000001";
			when "1111011111" => data_o <= "11111111000000000001";
			when "1111100000" => data_o <= "11111111000000000001";
			when "1111100001" => data_o <= "11111111000000000001";
			when "1111100010" => data_o <= "11111111000000000001";
			when "1111100011" => data_o <= "11111111000000000001";
			when "1111100100" => data_o <= "11111111000000000001";
			when "1111100101" => data_o <= "11111111000000000001";
			when "1111100110" => data_o <= "11111111000000000001";
			when "1111100111" => data_o <= "11111111000000000001";
			when "1111101000" => data_o <= "11111111000000000001";
			when "1111101001" => data_o <= "11111111000000000001";
			when "1111101010" => data_o <= "11111111000000000001";
			when "1111101011" => data_o <= "11111111000000000001";
			when "1111101100" => data_o <= "11111111000000000001";
			when "1111101101" => data_o <= "11111111000000000001";
			when "1111101110" => data_o <= "11111111000000000010";
			when "1111101111" => data_o <= "11111111000000000010";
			when "1111110000" => data_o <= "11111111000000000011";
			when "1111110001" => data_o <= "11111111000000000101";
			when "1111110010" => data_o <= "11111111000000001000";
			when "1111110011" => data_o <= "11111111000000001101";
			when "1111110100" => data_o <= "11111111000000010101";
			when "1111110101" => data_o <= "11111111000000100010";
			when "1111110110" => data_o <= "11111111000000110111";
			when "1111110111" => data_o <= "11111111000001011011";
			when "1111111000" => data_o <= "11111111000010010100";
			when "1111111001" => data_o <= "11111111000011110001";
			when "1111111010" => data_o <= "11111111000110000101";
			when "1111111011" => data_o <= "11111111001001101110";
			when "1111111100" => data_o <= "11111111001111010001";
			when "1111111101" => data_o <= "11111111010111010111";
			when "1111111110" => data_o <= "11111111100010011100";
			when "1111111111" => data_o <= "11111111110000010101";
			when "0000000000" => data_o <= "00000000000000000000";
			when "0000000001" => data_o <= "00000000001111101011";
			when "0000000010" => data_o <= "00000000011101100100";
			when "0000000011" => data_o <= "00000000101000101001";
			when "0000000100" => data_o <= "00000000110000101111";
			when "0000000101" => data_o <= "00000000110110010010";
			when "0000000110" => data_o <= "00000000111001111011";
			when "0000000111" => data_o <= "00000000111100001111";
			when "0000001000" => data_o <= "00000000111101101100";
			when "0000001001" => data_o <= "00000000111110100101";
			when "0000001010" => data_o <= "00000000111111001001";
			when "0000001011" => data_o <= "00000000111111011110";
			when "0000001100" => data_o <= "00000000111111101011";
			when "0000001101" => data_o <= "00000000111111110011";
			when "0000001110" => data_o <= "00000000111111111000";
			when "0000001111" => data_o <= "00000000111111111011";
			when "0000010000" => data_o <= "00000000111111111101";
			when "0000010001" => data_o <= "00000000111111111110";
			when "0000010010" => data_o <= "00000000111111111110";
			when "0000010011" => data_o <= "00000000111111111111";
			when "0000010100" => data_o <= "00000000111111111111";
			when "0000010101" => data_o <= "00000000111111111111";
			when "0000010110" => data_o <= "00000000111111111111";
			when "0000010111" => data_o <= "00000000111111111111";
			when "0000011000" => data_o <= "00000000111111111111";
			when "0000011001" => data_o <= "00000000111111111111";
			when "0000011010" => data_o <= "00000000111111111111";
			when "0000011011" => data_o <= "00000000111111111111";
			when "0000011100" => data_o <= "00000000111111111111";
			when "0000011101" => data_o <= "00000000111111111111";
			when "0000011110" => data_o <= "00000000111111111111";
			when "0000011111" => data_o <= "00000000111111111111";
			when "0000100000" => data_o <= "00000000111111111111";
			when "0000100001" => data_o <= "00000000111111111111";
			when "0000100010" => data_o <= "00000000111111111111";
			when "0000100011" => data_o <= "00000000111111111111";
			when "0000100100" => data_o <= "00000000111111111111";
			when "0000100101" => data_o <= "00000000111111111111";
			when "0000100110" => data_o <= "00000000111111111111";
			when "0000100111" => data_o <= "00000000111111111111";
			when "0000101000" => data_o <= "00000000111111111111";
			when "0000101001" => data_o <= "00000000111111111111";
			when "0000101010" => data_o <= "00000000111111111111";
			when "0000101011" => data_o <= "00000000111111111111";
			when "0000101100" => data_o <= "00000000111111111111";
			when "0000101101" => data_o <= "00000000111111111111";
			when "0000101110" => data_o <= "00000000111111111111";
			when "0000101111" => data_o <= "00000000111111111111";
			when "0000110000" => data_o <= "00000000111111111111";
			when "0000110001" => data_o <= "00000000111111111111";
			when "0000110010" => data_o <= "00000000111111111111";
			when "0000110011" => data_o <= "00000000111111111111";
			when "0000110100" => data_o <= "00000000111111111111";
			when "0000110101" => data_o <= "00000000111111111111";
			when "0000110110" => data_o <= "00000000111111111111";
			when "0000110111" => data_o <= "00000000111111111111";
			when "0000111000" => data_o <= "00000000111111111111";
			when "0000111001" => data_o <= "00000000111111111111";
			when "0000111010" => data_o <= "00000000111111111111";
			when "0000111011" => data_o <= "00000000111111111111";
			when "0000111100" => data_o <= "00000000111111111111";
			when "0000111101" => data_o <= "00000000111111111111";
			when "0000111110" => data_o <= "00000000111111111111";
			when "0000111111" => data_o <= "00000000111111111111";
			when "0001000000" => data_o <= "00000000111111111111";
			when "0001000001" => data_o <= "00000000111111111111";
			when "0001000010" => data_o <= "00000000111111111111";
			when "0001000011" => data_o <= "00000000111111111111";
			when "0001000100" => data_o <= "00000000111111111111";
			when "0001000101" => data_o <= "00000000111111111111";
			when "0001000110" => data_o <= "00000000111111111111";
			when "0001000111" => data_o <= "00000000111111111111";
			when "0001001000" => data_o <= "00000000111111111111";
			when "0001001001" => data_o <= "00000000111111111111";
			when "0001001010" => data_o <= "00000000111111111111";
			when "0001001011" => data_o <= "00000001000000000000";
			when "0001001100" => data_o <= "00000001000000000000";
			when "0001001101" => data_o <= "00000001000000000000";
			when "0001001110" => data_o <= "00000001000000000000";
			when "0001001111" => data_o <= "00000001000000000000";
			when "0001010000" => data_o <= "00000001000000000000";
			when "0001010001" => data_o <= "00000001000000000000";
			when "0001010010" => data_o <= "00000001000000000000";
			when "0001010011" => data_o <= "00000001000000000000";
			when "0001010100" => data_o <= "00000001000000000000";
			when "0001010101" => data_o <= "00000001000000000000";
			when "0001010110" => data_o <= "00000001000000000000";
			when "0001010111" => data_o <= "00000001000000000000";
			when "0001011000" => data_o <= "00000001000000000000";
			when "0001011001" => data_o <= "00000001000000000000";
			when "0001011010" => data_o <= "00000001000000000000";
			when "0001011011" => data_o <= "00000001000000000000";
			when "0001011100" => data_o <= "00000001000000000000";
			when "0001011101" => data_o <= "00000001000000000000";
			when "0001011110" => data_o <= "00000001000000000000";
			when "0001011111" => data_o <= "00000001000000000000";
			when "0001100000" => data_o <= "00000001000000000000";
			when "0001100001" => data_o <= "00000001000000000000";
			when "0001100010" => data_o <= "00000001000000000000";
			when "0001100011" => data_o <= "00000001000000000000";
			when "0001100100" => data_o <= "00000001000000000000";
			when "0001100101" => data_o <= "00000001000000000000";
			when "0001100110" => data_o <= "00000001000000000000";
			when "0001100111" => data_o <= "00000001000000000000";
			when "0001101000" => data_o <= "00000001000000000000";
			when "0001101001" => data_o <= "00000001000000000000";
			when "0001101010" => data_o <= "00000001000000000000";
			when "0001101011" => data_o <= "00000001000000000000";
			when "0001101100" => data_o <= "00000001000000000000";
			when "0001101101" => data_o <= "00000001000000000000";
			when "0001101110" => data_o <= "00000001000000000000";
			when "0001101111" => data_o <= "00000001000000000000";
			when "0001110000" => data_o <= "00000001000000000000";
			when "0001110001" => data_o <= "00000001000000000000";
			when "0001110010" => data_o <= "00000001000000000000";
			when "0001110011" => data_o <= "00000001000000000000";
			when "0001110100" => data_o <= "00000001000000000000";
			when "0001110101" => data_o <= "00000001000000000000";
			when "0001110110" => data_o <= "00000001000000000000";
			when "0001110111" => data_o <= "00000001000000000000";
			when "0001111000" => data_o <= "00000001000000000000";
			when "0001111001" => data_o <= "00000001000000000000";
			when "0001111010" => data_o <= "00000001000000000000";
			when "0001111011" => data_o <= "00000001000000000000";
			when "0001111100" => data_o <= "00000001000000000000";
			when "0001111101" => data_o <= "00000001000000000000";
			when "0001111110" => data_o <= "00000001000000000000";
			when "0001111111" => data_o <= "00000001000000000000";
			when "0010000000" => data_o <= "00000001000000000000";
			when "0010000001" => data_o <= "00000001000000000000";
			when "0010000010" => data_o <= "00000001000000000000";
			when "0010000011" => data_o <= "00000001000000000000";
			when "0010000100" => data_o <= "00000001000000000000";
			when "0010000101" => data_o <= "00000001000000000000";
			when "0010000110" => data_o <= "00000001000000000000";
			when "0010000111" => data_o <= "00000001000000000000";
			when "0010001000" => data_o <= "00000001000000000000";
			when "0010001001" => data_o <= "00000001000000000000";
			when "0010001010" => data_o <= "00000001000000000000";
			when "0010001011" => data_o <= "00000001000000000000";
			when "0010001100" => data_o <= "00000001000000000000";
			when "0010001101" => data_o <= "00000001000000000000";
			when "0010001110" => data_o <= "00000001000000000000";
			when "0010001111" => data_o <= "00000001000000000000";
			when "0010010000" => data_o <= "00000001000000000000";
			when "0010010001" => data_o <= "00000001000000000000";
			when "0010010010" => data_o <= "00000001000000000000";
			when "0010010011" => data_o <= "00000001000000000000";
			when "0010010100" => data_o <= "00000001000000000000";
			when "0010010101" => data_o <= "00000001000000000000";
			when "0010010110" => data_o <= "00000001000000000000";
			when "0010010111" => data_o <= "00000001000000000000";
			when "0010011000" => data_o <= "00000001000000000000";
			when "0010011001" => data_o <= "00000001000000000000";
			when "0010011010" => data_o <= "00000001000000000000";
			when "0010011011" => data_o <= "00000001000000000000";
			when "0010011100" => data_o <= "00000001000000000000";
			when "0010011101" => data_o <= "00000001000000000000";
			when "0010011110" => data_o <= "00000001000000000000";
			when "0010011111" => data_o <= "00000001000000000000";
			when "0010100000" => data_o <= "00000001000000000000";
			when "0010100001" => data_o <= "00000001000000000000";
			when "0010100010" => data_o <= "00000001000000000000";
			when "0010100011" => data_o <= "00000001000000000000";
			when "0010100100" => data_o <= "00000001000000000000";
			when "0010100101" => data_o <= "00000001000000000000";
			when "0010100110" => data_o <= "00000001000000000000";
			when "0010100111" => data_o <= "00000001000000000000";
			when "0010101000" => data_o <= "00000001000000000000";
			when "0010101001" => data_o <= "00000001000000000000";
			when "0010101010" => data_o <= "00000001000000000000";
			when "0010101011" => data_o <= "00000001000000000000";
			when "0010101100" => data_o <= "00000001000000000000";
			when "0010101101" => data_o <= "00000001000000000000";
			when "0010101110" => data_o <= "00000001000000000000";
			when "0010101111" => data_o <= "00000001000000000000";
			when "0010110000" => data_o <= "00000001000000000000";
			when "0010110001" => data_o <= "00000001000000000000";
			when "0010110010" => data_o <= "00000001000000000000";
			when "0010110011" => data_o <= "00000001000000000000";
			when "0010110100" => data_o <= "00000001000000000000";
			when "0010110101" => data_o <= "00000001000000000000";
			when "0010110110" => data_o <= "00000001000000000000";
			when "0010110111" => data_o <= "00000001000000000000";
			when "0010111000" => data_o <= "00000001000000000000";
			when "0010111001" => data_o <= "00000001000000000000";
			when "0010111010" => data_o <= "00000001000000000000";
			when "0010111011" => data_o <= "00000001000000000000";
			when "0010111100" => data_o <= "00000001000000000000";
			when "0010111101" => data_o <= "00000001000000000000";
			when "0010111110" => data_o <= "00000001000000000000";
			when "0010111111" => data_o <= "00000001000000000000";
			when "0011000000" => data_o <= "00000001000000000000";
			when "0011000001" => data_o <= "00000001000000000000";
			when "0011000010" => data_o <= "00000001000000000000";
			when "0011000011" => data_o <= "00000001000000000000";
			when "0011000100" => data_o <= "00000001000000000000";
			when "0011000101" => data_o <= "00000001000000000000";
			when "0011000110" => data_o <= "00000001000000000000";
			when "0011000111" => data_o <= "00000001000000000000";
			when "0011001000" => data_o <= "00000001000000000000";
			when "0011001001" => data_o <= "00000001000000000000";
			when "0011001010" => data_o <= "00000001000000000000";
			when "0011001011" => data_o <= "00000001000000000000";
			when "0011001100" => data_o <= "00000001000000000000";
			when "0011001101" => data_o <= "00000001000000000000";
			when "0011001110" => data_o <= "00000001000000000000";
			when "0011001111" => data_o <= "00000001000000000000";
			when "0011010000" => data_o <= "00000001000000000000";
			when "0011010001" => data_o <= "00000001000000000000";
			when "0011010010" => data_o <= "00000001000000000000";
			when "0011010011" => data_o <= "00000001000000000000";
			when "0011010100" => data_o <= "00000001000000000000";
			when "0011010101" => data_o <= "00000001000000000000";
			when "0011010110" => data_o <= "00000001000000000000";
			when "0011010111" => data_o <= "00000001000000000000";
			when "0011011000" => data_o <= "00000001000000000000";
			when "0011011001" => data_o <= "00000001000000000000";
			when "0011011010" => data_o <= "00000001000000000000";
			when "0011011011" => data_o <= "00000001000000000000";
			when "0011011100" => data_o <= "00000001000000000000";
			when "0011011101" => data_o <= "00000001000000000000";
			when "0011011110" => data_o <= "00000001000000000000";
			when "0011011111" => data_o <= "00000001000000000000";
			when "0011100000" => data_o <= "00000001000000000000";
			when "0011100001" => data_o <= "00000001000000000000";
			when "0011100010" => data_o <= "00000001000000000000";
			when "0011100011" => data_o <= "00000001000000000000";
			when "0011100100" => data_o <= "00000001000000000000";
			when "0011100101" => data_o <= "00000001000000000000";
			when "0011100110" => data_o <= "00000001000000000000";
			when "0011100111" => data_o <= "00000001000000000000";
			when "0011101000" => data_o <= "00000001000000000000";
			when "0011101001" => data_o <= "00000001000000000000";
			when "0011101010" => data_o <= "00000001000000000000";
			when "0011101011" => data_o <= "00000001000000000000";
			when "0011101100" => data_o <= "00000001000000000000";
			when "0011101101" => data_o <= "00000001000000000000";
			when "0011101110" => data_o <= "00000001000000000000";
			when "0011101111" => data_o <= "00000001000000000000";
			when "0011110000" => data_o <= "00000001000000000000";
			when "0011110001" => data_o <= "00000001000000000000";
			when "0011110010" => data_o <= "00000001000000000000";
			when "0011110011" => data_o <= "00000001000000000000";
			when "0011110100" => data_o <= "00000001000000000000";
			when "0011110101" => data_o <= "00000001000000000000";
			when "0011110110" => data_o <= "00000001000000000000";
			when "0011110111" => data_o <= "00000001000000000000";
			when "0011111000" => data_o <= "00000001000000000000";
			when "0011111001" => data_o <= "00000001000000000000";
			when "0011111010" => data_o <= "00000001000000000000";
			when "0011111011" => data_o <= "00000001000000000000";
			when "0011111100" => data_o <= "00000001000000000000";
			when "0011111101" => data_o <= "00000001000000000000";
			when "0011111110" => data_o <= "00000001000000000000";
			when "0011111111" => data_o <= "00000001000000000000";
			when "0100000000" => data_o <= "00000001000000000000";
			when "0100000001" => data_o <= "00000001000000000000";
			when "0100000010" => data_o <= "00000001000000000000";
			when "0100000011" => data_o <= "00000001000000000000";
			when "0100000100" => data_o <= "00000001000000000000";
			when "0100000101" => data_o <= "00000001000000000000";
			when "0100000110" => data_o <= "00000001000000000000";
			when "0100000111" => data_o <= "00000001000000000000";
			when "0100001000" => data_o <= "00000001000000000000";
			when "0100001001" => data_o <= "00000001000000000000";
			when "0100001010" => data_o <= "00000001000000000000";
			when "0100001011" => data_o <= "00000001000000000000";
			when "0100001100" => data_o <= "00000001000000000000";
			when "0100001101" => data_o <= "00000001000000000000";
			when "0100001110" => data_o <= "00000001000000000000";
			when "0100001111" => data_o <= "00000001000000000000";
			when "0100010000" => data_o <= "00000001000000000000";
			when "0100010001" => data_o <= "00000001000000000000";
			when "0100010010" => data_o <= "00000001000000000000";
			when "0100010011" => data_o <= "00000001000000000000";
			when "0100010100" => data_o <= "00000001000000000000";
			when "0100010101" => data_o <= "00000001000000000000";
			when "0100010110" => data_o <= "00000001000000000000";
			when "0100010111" => data_o <= "00000001000000000000";
			when "0100011000" => data_o <= "00000001000000000000";
			when "0100011001" => data_o <= "00000001000000000000";
			when "0100011010" => data_o <= "00000001000000000000";
			when "0100011011" => data_o <= "00000001000000000000";
			when "0100011100" => data_o <= "00000001000000000000";
			when "0100011101" => data_o <= "00000001000000000000";
			when "0100011110" => data_o <= "00000001000000000000";
			when "0100011111" => data_o <= "00000001000000000000";
			when "0100100000" => data_o <= "00000001000000000000";
			when "0100100001" => data_o <= "00000001000000000000";
			when "0100100010" => data_o <= "00000001000000000000";
			when "0100100011" => data_o <= "00000001000000000000";
			when "0100100100" => data_o <= "00000001000000000000";
			when "0100100101" => data_o <= "00000001000000000000";
			when "0100100110" => data_o <= "00000001000000000000";
			when "0100100111" => data_o <= "00000001000000000000";
			when "0100101000" => data_o <= "00000001000000000000";
			when "0100101001" => data_o <= "00000001000000000000";
			when "0100101010" => data_o <= "00000001000000000000";
			when "0100101011" => data_o <= "00000001000000000000";
			when "0100101100" => data_o <= "00000001000000000000";
			when "0100101101" => data_o <= "00000001000000000000";
			when "0100101110" => data_o <= "00000001000000000000";
			when "0100101111" => data_o <= "00000001000000000000";
			when "0100110000" => data_o <= "00000001000000000000";
			when "0100110001" => data_o <= "00000001000000000000";
			when "0100110010" => data_o <= "00000001000000000000";
			when "0100110011" => data_o <= "00000001000000000000";
			when "0100110100" => data_o <= "00000001000000000000";
			when "0100110101" => data_o <= "00000001000000000000";
			when "0100110110" => data_o <= "00000001000000000000";
			when "0100110111" => data_o <= "00000001000000000000";
			when "0100111000" => data_o <= "00000001000000000000";
			when "0100111001" => data_o <= "00000001000000000000";
			when "0100111010" => data_o <= "00000001000000000000";
			when "0100111011" => data_o <= "00000001000000000000";
			when "0100111100" => data_o <= "00000001000000000000";
			when "0100111101" => data_o <= "00000001000000000000";
			when "0100111110" => data_o <= "00000001000000000000";
			when "0100111111" => data_o <= "00000001000000000000";
			when "0101000000" => data_o <= "00000001000000000000";
			when "0101000001" => data_o <= "00000001000000000000";
			when "0101000010" => data_o <= "00000001000000000000";
			when "0101000011" => data_o <= "00000001000000000000";
			when "0101000100" => data_o <= "00000001000000000000";
			when "0101000101" => data_o <= "00000001000000000000";
			when "0101000110" => data_o <= "00000001000000000000";
			when "0101000111" => data_o <= "00000001000000000000";
			when "0101001000" => data_o <= "00000001000000000000";
			when "0101001001" => data_o <= "00000001000000000000";
			when "0101001010" => data_o <= "00000001000000000000";
			when "0101001011" => data_o <= "00000001000000000000";
			when "0101001100" => data_o <= "00000001000000000000";
			when "0101001101" => data_o <= "00000001000000000000";
			when "0101001110" => data_o <= "00000001000000000000";
			when "0101001111" => data_o <= "00000001000000000000";
			when "0101010000" => data_o <= "00000001000000000000";
			when "0101010001" => data_o <= "00000001000000000000";
			when "0101010010" => data_o <= "00000001000000000000";
			when "0101010011" => data_o <= "00000001000000000000";
			when "0101010100" => data_o <= "00000001000000000000";
			when "0101010101" => data_o <= "00000001000000000000";
			when "0101010110" => data_o <= "00000001000000000000";
			when "0101010111" => data_o <= "00000001000000000000";
			when "0101011000" => data_o <= "00000001000000000000";
			when "0101011001" => data_o <= "00000001000000000000";
			when "0101011010" => data_o <= "00000001000000000000";
			when "0101011011" => data_o <= "00000001000000000000";
			when "0101011100" => data_o <= "00000001000000000000";
			when "0101011101" => data_o <= "00000001000000000000";
			when "0101011110" => data_o <= "00000001000000000000";
			when "0101011111" => data_o <= "00000001000000000000";
			when "0101100000" => data_o <= "00000001000000000000";
			when "0101100001" => data_o <= "00000001000000000000";
			when "0101100010" => data_o <= "00000001000000000000";
			when "0101100011" => data_o <= "00000001000000000000";
			when "0101100100" => data_o <= "00000001000000000000";
			when "0101100101" => data_o <= "00000001000000000000";
			when "0101100110" => data_o <= "00000001000000000000";
			when "0101100111" => data_o <= "00000001000000000000";
			when "0101101000" => data_o <= "00000001000000000000";
			when "0101101001" => data_o <= "00000001000000000000";
			when "0101101010" => data_o <= "00000001000000000000";
			when "0101101011" => data_o <= "00000001000000000000";
			when "0101101100" => data_o <= "00000001000000000000";
			when "0101101101" => data_o <= "00000001000000000000";
			when "0101101110" => data_o <= "00000001000000000000";
			when "0101101111" => data_o <= "00000001000000000000";
			when "0101110000" => data_o <= "00000001000000000000";
			when "0101110001" => data_o <= "00000001000000000000";
			when "0101110010" => data_o <= "00000001000000000000";
			when "0101110011" => data_o <= "00000001000000000000";
			when "0101110100" => data_o <= "00000001000000000000";
			when "0101110101" => data_o <= "00000001000000000000";
			when "0101110110" => data_o <= "00000001000000000000";
			when "0101110111" => data_o <= "00000001000000000000";
			when "0101111000" => data_o <= "00000001000000000000";
			when "0101111001" => data_o <= "00000001000000000000";
			when "0101111010" => data_o <= "00000001000000000000";
			when "0101111011" => data_o <= "00000001000000000000";
			when "0101111100" => data_o <= "00000001000000000000";
			when "0101111101" => data_o <= "00000001000000000000";
			when "0101111110" => data_o <= "00000001000000000000";
			when "0101111111" => data_o <= "00000001000000000000";
			when "0110000000" => data_o <= "00000001000000000000";
			when "0110000001" => data_o <= "00000001000000000000";
			when "0110000010" => data_o <= "00000001000000000000";
			when "0110000011" => data_o <= "00000001000000000000";
			when "0110000100" => data_o <= "00000001000000000000";
			when "0110000101" => data_o <= "00000001000000000000";
			when "0110000110" => data_o <= "00000001000000000000";
			when "0110000111" => data_o <= "00000001000000000000";
			when "0110001000" => data_o <= "00000001000000000000";
			when "0110001001" => data_o <= "00000001000000000000";
			when "0110001010" => data_o <= "00000001000000000000";
			when "0110001011" => data_o <= "00000001000000000000";
			when "0110001100" => data_o <= "00000001000000000000";
			when "0110001101" => data_o <= "00000001000000000000";
			when "0110001110" => data_o <= "00000001000000000000";
			when "0110001111" => data_o <= "00000001000000000000";
			when "0110010000" => data_o <= "00000001000000000000";
			when "0110010001" => data_o <= "00000001000000000000";
			when "0110010010" => data_o <= "00000001000000000000";
			when "0110010011" => data_o <= "00000001000000000000";
			when "0110010100" => data_o <= "00000001000000000000";
			when "0110010101" => data_o <= "00000001000000000000";
			when "0110010110" => data_o <= "00000001000000000000";
			when "0110010111" => data_o <= "00000001000000000000";
			when "0110011000" => data_o <= "00000001000000000000";
			when "0110011001" => data_o <= "00000001000000000000";
			when "0110011010" => data_o <= "00000001000000000000";
			when "0110011011" => data_o <= "00000001000000000000";
			when "0110011100" => data_o <= "00000001000000000000";
			when "0110011101" => data_o <= "00000001000000000000";
			when "0110011110" => data_o <= "00000001000000000000";
			when "0110011111" => data_o <= "00000001000000000000";
			when "0110100000" => data_o <= "00000001000000000000";
			when "0110100001" => data_o <= "00000001000000000000";
			when "0110100010" => data_o <= "00000001000000000000";
			when "0110100011" => data_o <= "00000001000000000000";
			when "0110100100" => data_o <= "00000001000000000000";
			when "0110100101" => data_o <= "00000001000000000000";
			when "0110100110" => data_o <= "00000001000000000000";
			when "0110100111" => data_o <= "00000001000000000000";
			when "0110101000" => data_o <= "00000001000000000000";
			when "0110101001" => data_o <= "00000001000000000000";
			when "0110101010" => data_o <= "00000001000000000000";
			when "0110101011" => data_o <= "00000001000000000000";
			when "0110101100" => data_o <= "00000001000000000000";
			when "0110101101" => data_o <= "00000001000000000000";
			when "0110101110" => data_o <= "00000001000000000000";
			when "0110101111" => data_o <= "00000001000000000000";
			when "0110110000" => data_o <= "00000001000000000000";
			when "0110110001" => data_o <= "00000001000000000000";
			when "0110110010" => data_o <= "00000001000000000000";
			when "0110110011" => data_o <= "00000001000000000000";
			when "0110110100" => data_o <= "00000001000000000000";
			when "0110110101" => data_o <= "00000001000000000000";
			when "0110110110" => data_o <= "00000001000000000000";
			when "0110110111" => data_o <= "00000001000000000000";
			when "0110111000" => data_o <= "00000001000000000000";
			when "0110111001" => data_o <= "00000001000000000000";
			when "0110111010" => data_o <= "00000001000000000000";
			when "0110111011" => data_o <= "00000001000000000000";
			when "0110111100" => data_o <= "00000001000000000000";
			when "0110111101" => data_o <= "00000001000000000000";
			when "0110111110" => data_o <= "00000001000000000000";
			when "0110111111" => data_o <= "00000001000000000000";
			when "0111000000" => data_o <= "00000001000000000000";
			when "0111000001" => data_o <= "00000001000000000000";
			when "0111000010" => data_o <= "00000001000000000000";
			when "0111000011" => data_o <= "00000001000000000000";
			when "0111000100" => data_o <= "00000001000000000000";
			when "0111000101" => data_o <= "00000001000000000000";
			when "0111000110" => data_o <= "00000001000000000000";
			when "0111000111" => data_o <= "00000001000000000000";
			when "0111001000" => data_o <= "00000001000000000000";
			when "0111001001" => data_o <= "00000001000000000000";
			when "0111001010" => data_o <= "00000001000000000000";
			when "0111001011" => data_o <= "00000001000000000000";
			when "0111001100" => data_o <= "00000001000000000000";
			when "0111001101" => data_o <= "00000001000000000000";
			when "0111001110" => data_o <= "00000001000000000000";
			when "0111001111" => data_o <= "00000001000000000000";
			when "0111010000" => data_o <= "00000001000000000000";
			when "0111010001" => data_o <= "00000001000000000000";
			when "0111010010" => data_o <= "00000001000000000000";
			when "0111010011" => data_o <= "00000001000000000000";
			when "0111010100" => data_o <= "00000001000000000000";
			when "0111010101" => data_o <= "00000001000000000000";
			when "0111010110" => data_o <= "00000001000000000000";
			when "0111010111" => data_o <= "00000001000000000000";
			when "0111011000" => data_o <= "00000001000000000000";
			when "0111011001" => data_o <= "00000001000000000000";
			when "0111011010" => data_o <= "00000001000000000000";
			when "0111011011" => data_o <= "00000001000000000000";
			when "0111011100" => data_o <= "00000001000000000000";
			when "0111011101" => data_o <= "00000001000000000000";
			when "0111011110" => data_o <= "00000001000000000000";
			when "0111011111" => data_o <= "00000001000000000000";
			when "0111100000" => data_o <= "00000001000000000000";
			when "0111100001" => data_o <= "00000001000000000000";
			when "0111100010" => data_o <= "00000001000000000000";
			when "0111100011" => data_o <= "00000001000000000000";
			when "0111100100" => data_o <= "00000001000000000000";
			when "0111100101" => data_o <= "00000001000000000000";
			when "0111100110" => data_o <= "00000001000000000000";
			when "0111100111" => data_o <= "00000001000000000000";
			when "0111101000" => data_o <= "00000001000000000000";
			when "0111101001" => data_o <= "00000001000000000000";
			when "0111101010" => data_o <= "00000001000000000000";
			when "0111101011" => data_o <= "00000001000000000000";
			when "0111101100" => data_o <= "00000001000000000000";
			when "0111101101" => data_o <= "00000001000000000000";
			when "0111101110" => data_o <= "00000001000000000000";
			when "0111101111" => data_o <= "00000001000000000000";
			when "0111110000" => data_o <= "00000001000000000000";
			when "0111110001" => data_o <= "00000001000000000000";
			when "0111110010" => data_o <= "00000001000000000000";
			when "0111110011" => data_o <= "00000001000000000000";
			when "0111110100" => data_o <= "00000001000000000000";
			when "0111110101" => data_o <= "00000001000000000000";
			when "0111110110" => data_o <= "00000001000000000000";
			when "0111110111" => data_o <= "00000001000000000000";
			when "0111111000" => data_o <= "00000001000000000000";
			when "0111111001" => data_o <= "00000001000000000000";
			when "0111111010" => data_o <= "00000001000000000000";
			when "0111111011" => data_o <= "00000001000000000000";
			when "0111111100" => data_o <= "00000001000000000000";
			when "0111111101" => data_o <= "00000001000000000000";
			when "0111111110" => data_o <= "00000001000000000000";
			when "0111111111" => data_o <= "00000001000000000000";
			when others => data_o <= "00000000000000000000";
		end case;
	end process;
end architecture;
